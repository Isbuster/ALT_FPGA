-- my_MCU.vhd

-- Generated using ACDS version 23.1 993

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity my_MCU is
	port (
		clk_clk            : in    std_logic                     := '0';             --         clk.clk
		i2c_scl            : out   std_logic;                                        --         i2c.scl
		i2c_sda            : inout std_logic                     := '0';             --            .sda
		pio_in_ext_export  : in    std_logic_vector(15 downto 0) := (others => '0'); --  pio_in_ext.export
		pio_out_ext_export : out   std_logic_vector(15 downto 0);                    -- pio_out_ext.export
		reset_reset_n      : in    std_logic                     := '0'              --       reset.reset_n
	);
end entity my_MCU;

architecture rtl of my_MCU is
	component I2C_MASTER_ALL is
		port (
			CLK        : in    std_logic                     := 'X';             -- clk
			chipselect : in    std_logic                     := 'X';             -- chipselect
			wr         : in    std_logic                     := 'X';             -- write
			rd         : in    std_logic                     := 'X';             -- read
			address    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			scl        : out   std_logic;                                        -- scl
			sda        : inout std_logic                     := 'X';             -- sda
			RST        : in    std_logic                     := 'X'              -- reset
		);
	end component I2C_MASTER_ALL;

	component my_MCU_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component my_MCU_jtag;

	component my_MCU_nios is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component my_MCU_nios;

	component my_MCU_pio_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component my_MCU_pio_in;

	component my_MCU_pio_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component my_MCU_pio_out;

	component my_MCU_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component my_MCU_ram;

	component my_MCU_mm_interconnect_0 is
		port (
			clk_0_clk_clk                          : in  std_logic                     := 'X';             -- clk
			nios_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios_data_master_address               : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			nios_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios_instruction_master_address        : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			nios_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			I2C_MASTER_5_avalon_slave_0_address    : out std_logic_vector(2 downto 0);                     -- address
			I2C_MASTER_5_avalon_slave_0_write      : out std_logic;                                        -- write
			I2C_MASTER_5_avalon_slave_0_read       : out std_logic;                                        -- read
			I2C_MASTER_5_avalon_slave_0_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			I2C_MASTER_5_avalon_slave_0_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			I2C_MASTER_5_avalon_slave_0_chipselect : out std_logic;                                        -- chipselect
			jtag_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			nios_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios_debug_mem_slave_write             : out std_logic;                                        -- write
			nios_debug_mem_slave_read              : out std_logic;                                        -- read
			nios_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			pio_in_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			pio_in_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			pio_out_s1_write                       : out std_logic;                                        -- write
			pio_out_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_out_s1_chipselect                  : out std_logic;                                        -- chipselect
			ram_s1_address                         : out std_logic_vector(15 downto 0);                    -- address
			ram_s1_write                           : out std_logic;                                        -- write
			ram_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ram_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			ram_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			ram_s1_chipselect                      : out std_logic;                                        -- chipselect
			ram_s1_clken                           : out std_logic                                         -- clken
		);
	end component my_MCU_mm_interconnect_0;

	component my_MCU_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component my_MCU_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios_data_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	signal nios_data_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	signal nios_data_master_debugaccess                             : std_logic;                     -- nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	signal nios_data_master_address                                 : std_logic_vector(19 downto 0); -- nios:d_address -> mm_interconnect_0:nios_data_master_address
	signal nios_data_master_byteenable                              : std_logic_vector(3 downto 0);  -- nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	signal nios_data_master_read                                    : std_logic;                     -- nios:d_read -> mm_interconnect_0:nios_data_master_read
	signal nios_data_master_write                                   : std_logic;                     -- nios:d_write -> mm_interconnect_0:nios_data_master_write
	signal nios_data_master_writedata                               : std_logic_vector(31 downto 0); -- nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	signal nios_instruction_master_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	signal nios_instruction_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	signal nios_instruction_master_address                          : std_logic_vector(19 downto 0); -- nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	signal nios_instruction_master_read                             : std_logic;                     -- nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	signal mm_interconnect_0_i2c_master_5_avalon_slave_0_chipselect : std_logic;                     -- mm_interconnect_0:I2C_MASTER_5_avalon_slave_0_chipselect -> I2C_MASTER_5:chipselect
	signal mm_interconnect_0_i2c_master_5_avalon_slave_0_readdata   : std_logic_vector(31 downto 0); -- I2C_MASTER_5:readdata -> mm_interconnect_0:I2C_MASTER_5_avalon_slave_0_readdata
	signal mm_interconnect_0_i2c_master_5_avalon_slave_0_address    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:I2C_MASTER_5_avalon_slave_0_address -> I2C_MASTER_5:address
	signal mm_interconnect_0_i2c_master_5_avalon_slave_0_read       : std_logic;                     -- mm_interconnect_0:I2C_MASTER_5_avalon_slave_0_read -> I2C_MASTER_5:rd
	signal mm_interconnect_0_i2c_master_5_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:I2C_MASTER_5_avalon_slave_0_write -> I2C_MASTER_5:wr
	signal mm_interconnect_0_i2c_master_5_avalon_slave_0_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:I2C_MASTER_5_avalon_slave_0_writedata -> I2C_MASTER_5:writedata
	signal mm_interconnect_0_nios_debug_mem_slave_readdata          : std_logic_vector(31 downto 0); -- nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_debug_mem_slave_waitrequest       : std_logic;                     -- nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_debug_mem_slave_debugaccess       : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_debug_mem_slave_address           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	signal mm_interconnect_0_nios_debug_mem_slave_read              : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	signal mm_interconnect_0_nios_debug_mem_slave_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_debug_mem_slave_write             : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	signal mm_interconnect_0_nios_debug_mem_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	signal mm_interconnect_0_ram_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	signal mm_interconnect_0_ram_s1_readdata                        : std_logic_vector(31 downto 0); -- ram:readdata -> mm_interconnect_0:ram_s1_readdata
	signal mm_interconnect_0_ram_s1_address                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:ram_s1_address -> ram:address
	signal mm_interconnect_0_ram_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	signal mm_interconnect_0_ram_s1_write                           : std_logic;                     -- mm_interconnect_0:ram_s1_write -> ram:write
	signal mm_interconnect_0_ram_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:ram_s1_writedata -> ram:writedata
	signal mm_interconnect_0_ram_s1_clken                           : std_logic;                     -- mm_interconnect_0:ram_s1_clken -> ram:clken
	signal mm_interconnect_0_pio_in_s1_readdata                     : std_logic_vector(31 downto 0); -- pio_in:readdata -> mm_interconnect_0:pio_in_s1_readdata
	signal mm_interconnect_0_pio_in_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_in_s1_address -> pio_in:address
	signal mm_interconnect_0_pio_out_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:pio_out_s1_chipselect -> pio_out:chipselect
	signal mm_interconnect_0_pio_out_s1_readdata                    : std_logic_vector(31 downto 0); -- pio_out:readdata -> mm_interconnect_0:pio_out_s1_readdata
	signal mm_interconnect_0_pio_out_s1_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_out_s1_address -> pio_out:address
	signal mm_interconnect_0_pio_out_s1_write                       : std_logic;                     -- mm_interconnect_0:pio_out_s1_write -> mm_interconnect_0_pio_out_s1_write:in
	signal mm_interconnect_0_pio_out_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_out_s1_writedata -> pio_out:writedata
	signal irq_mapper_receiver0_irq                                 : std_logic;                     -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal nios_irq_irq                                             : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios:irq
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [I2C_MASTER_5:RST, irq_mapper:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                       : std_logic;                     -- rst_controller:reset_req -> [nios:reset_req, ram:reset_req, rst_translator:reset_req_in]
	signal nios_debug_reset_request_reset                           : std_logic;                     -- nios:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                  : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> jtag:av_read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> jtag:av_write_n
	signal mm_interconnect_0_pio_out_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_pio_out_s1_write:inv -> pio_out:write_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag:rst_n, nios:reset_n, pio_in:reset_n, pio_out:reset_n]

begin

	i2c_master_5 : component I2C_MASTER_ALL
		port map (
			CLK        => clk_clk,                                                  --          clock.clk
			chipselect => mm_interconnect_0_i2c_master_5_avalon_slave_0_chipselect, -- avalon_slave_0.chipselect
			wr         => mm_interconnect_0_i2c_master_5_avalon_slave_0_write,      --               .write
			rd         => mm_interconnect_0_i2c_master_5_avalon_slave_0_read,       --               .read
			address    => mm_interconnect_0_i2c_master_5_avalon_slave_0_address,    --               .address
			writedata  => mm_interconnect_0_i2c_master_5_avalon_slave_0_writedata,  --               .writedata
			readdata   => mm_interconnect_0_i2c_master_5_avalon_slave_0_readdata,   --               .readdata
			scl        => i2c_scl,                                                  --    conduit_end.scl
			sda        => i2c_sda,                                                  --               .sda
			RST        => rst_controller_reset_out_reset                            --     reset_sink.reset
		);

	jtag : component my_MCU_jtag
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	nios : component my_MCU_nios
		port map (
			clk                                 => clk_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,           --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                 --                          .reset_req
			d_address                           => nios_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_data_master_read,                              --                          .read
			d_readdata                          => nios_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_data_master_write,                             --                          .write
			d_writedata                         => nios_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_instruction_master_read,                       --                          .read
			i_readdata                          => nios_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                -- custom_instruction_master.readra
		);

	pio_in : component my_MCU_pio_in
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pio_in_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_pio_in_s1_readdata,     --                    .readdata
			in_port  => pio_in_ext_export                         -- external_connection.export
		);

	pio_out : component my_MCU_pio_out
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_out_s1_readdata,        --                    .readdata
			out_port   => pio_out_ext_export                            -- external_connection.export
		);

	ram : component my_MCU_ram
		port map (
			clk        => clk_clk,                             --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,  --       .reset_req
			freeze     => '0'                                  -- (terminated)
		);

	mm_interconnect_0 : component my_MCU_mm_interconnect_0
		port map (
			clk_0_clk_clk                          => clk_clk,                                                  --                        clk_0_clk.clk
			nios_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                           -- nios_reset_reset_bridge_in_reset.reset
			nios_data_master_address               => nios_data_master_address,                                 --                 nios_data_master.address
			nios_data_master_waitrequest           => nios_data_master_waitrequest,                             --                                 .waitrequest
			nios_data_master_byteenable            => nios_data_master_byteenable,                              --                                 .byteenable
			nios_data_master_read                  => nios_data_master_read,                                    --                                 .read
			nios_data_master_readdata              => nios_data_master_readdata,                                --                                 .readdata
			nios_data_master_write                 => nios_data_master_write,                                   --                                 .write
			nios_data_master_writedata             => nios_data_master_writedata,                               --                                 .writedata
			nios_data_master_debugaccess           => nios_data_master_debugaccess,                             --                                 .debugaccess
			nios_instruction_master_address        => nios_instruction_master_address,                          --          nios_instruction_master.address
			nios_instruction_master_waitrequest    => nios_instruction_master_waitrequest,                      --                                 .waitrequest
			nios_instruction_master_read           => nios_instruction_master_read,                             --                                 .read
			nios_instruction_master_readdata       => nios_instruction_master_readdata,                         --                                 .readdata
			I2C_MASTER_5_avalon_slave_0_address    => mm_interconnect_0_i2c_master_5_avalon_slave_0_address,    --      I2C_MASTER_5_avalon_slave_0.address
			I2C_MASTER_5_avalon_slave_0_write      => mm_interconnect_0_i2c_master_5_avalon_slave_0_write,      --                                 .write
			I2C_MASTER_5_avalon_slave_0_read       => mm_interconnect_0_i2c_master_5_avalon_slave_0_read,       --                                 .read
			I2C_MASTER_5_avalon_slave_0_readdata   => mm_interconnect_0_i2c_master_5_avalon_slave_0_readdata,   --                                 .readdata
			I2C_MASTER_5_avalon_slave_0_writedata  => mm_interconnect_0_i2c_master_5_avalon_slave_0_writedata,  --                                 .writedata
			I2C_MASTER_5_avalon_slave_0_chipselect => mm_interconnect_0_i2c_master_5_avalon_slave_0_chipselect, --                                 .chipselect
			jtag_avalon_jtag_slave_address         => mm_interconnect_0_jtag_avalon_jtag_slave_address,         --           jtag_avalon_jtag_slave.address
			jtag_avalon_jtag_slave_write           => mm_interconnect_0_jtag_avalon_jtag_slave_write,           --                                 .write
			jtag_avalon_jtag_slave_read            => mm_interconnect_0_jtag_avalon_jtag_slave_read,            --                                 .read
			jtag_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                                 .readdata
			jtag_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                                 .writedata
			jtag_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                                 .waitrequest
			jtag_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      --                                 .chipselect
			nios_debug_mem_slave_address           => mm_interconnect_0_nios_debug_mem_slave_address,           --             nios_debug_mem_slave.address
			nios_debug_mem_slave_write             => mm_interconnect_0_nios_debug_mem_slave_write,             --                                 .write
			nios_debug_mem_slave_read              => mm_interconnect_0_nios_debug_mem_slave_read,              --                                 .read
			nios_debug_mem_slave_readdata          => mm_interconnect_0_nios_debug_mem_slave_readdata,          --                                 .readdata
			nios_debug_mem_slave_writedata         => mm_interconnect_0_nios_debug_mem_slave_writedata,         --                                 .writedata
			nios_debug_mem_slave_byteenable        => mm_interconnect_0_nios_debug_mem_slave_byteenable,        --                                 .byteenable
			nios_debug_mem_slave_waitrequest       => mm_interconnect_0_nios_debug_mem_slave_waitrequest,       --                                 .waitrequest
			nios_debug_mem_slave_debugaccess       => mm_interconnect_0_nios_debug_mem_slave_debugaccess,       --                                 .debugaccess
			pio_in_s1_address                      => mm_interconnect_0_pio_in_s1_address,                      --                        pio_in_s1.address
			pio_in_s1_readdata                     => mm_interconnect_0_pio_in_s1_readdata,                     --                                 .readdata
			pio_out_s1_address                     => mm_interconnect_0_pio_out_s1_address,                     --                       pio_out_s1.address
			pio_out_s1_write                       => mm_interconnect_0_pio_out_s1_write,                       --                                 .write
			pio_out_s1_readdata                    => mm_interconnect_0_pio_out_s1_readdata,                    --                                 .readdata
			pio_out_s1_writedata                   => mm_interconnect_0_pio_out_s1_writedata,                   --                                 .writedata
			pio_out_s1_chipselect                  => mm_interconnect_0_pio_out_s1_chipselect,                  --                                 .chipselect
			ram_s1_address                         => mm_interconnect_0_ram_s1_address,                         --                           ram_s1.address
			ram_s1_write                           => mm_interconnect_0_ram_s1_write,                           --                                 .write
			ram_s1_readdata                        => mm_interconnect_0_ram_s1_readdata,                        --                                 .readdata
			ram_s1_writedata                       => mm_interconnect_0_ram_s1_writedata,                       --                                 .writedata
			ram_s1_byteenable                      => mm_interconnect_0_ram_s1_byteenable,                      --                                 .byteenable
			ram_s1_chipselect                      => mm_interconnect_0_ram_s1_chipselect,                      --                                 .chipselect
			ram_s1_clken                           => mm_interconnect_0_ram_s1_clken                            --                                 .clken
		);

	irq_mapper : component my_MCU_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios_irq_irq                    --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios_debug_reset_request_reset,     -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_pio_out_s1_write_ports_inv <= not mm_interconnect_0_pio_out_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of my_MCU
