pixel_clk_inst : pixel_clk PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
