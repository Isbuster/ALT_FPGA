LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

--GJELDER 60HZ 640x480
--
-- Pixel clock (MHz) = 25.175
--
-- Horizontal
-- Sync pulse = 96
-- Front porch = 16
-- Back porch = 48
-- Hsync polarity = n
-- 
-- Vertical 
-- Sync pulse = 2
-- Front porch = 10
-- Back porch = 33
-- Vsync polarity = n

ENTITY vga_testbrett IS
  PORT ( 
    clk         : IN STD_LOGIC;
    KEY         : IN STD_LOGIC_VECTOR(3 downto 0);
    VGA_CLK     : OUT STD_LOGIC;
    VGA_BLANK_N : OUT STD_LOGIC;
    VGA_SYNC_N  : OUT STD_LOGIC;
    VGA_HS      : OUT STD_LOGIC;
    VGA_VS      : OUT STD_LOGIC;
    VGA_R       : OUT STD_LOGIC_VECTOR(7 downto 0);
    VGA_G       : OUT STD_LOGIC_VECTOR(7 downto 0);
    VGA_B       : OUT STD_LOGIC_VECTOR(7 downto 0)
  );
END ENTITY;

ARCHITECTURE RTL OF vga_testbrett IS
  SIGNAL display_en : STD_LOGIC;
  SIGNAL column     : INTEGER;
  SIGNAL row        : INTEGER;

  COMPONENT vga_adapter IS
    PORT ( 
      pixel_clk   : IN  STD_LOGIC;
      reset_n     : IN  STD_LOGIC;
      h_sync      : OUT STD_LOGIC;
      v_sync      : OUT STD_LOGIC;
      blank_n     : OUT STD_LOGIC;
      sync_n      : OUT STD_LOGIC;
      display_en  : OUT STD_LOGIC;
      column      : OUT INTEGER;
      row         : OUT INTEGER
    );
  END COMPONENT;
BEGIN
  VGA_CLK <= clk;
  
  vga_square_test : process(display_en, row, column) is
    variable y_length : integer range 0 to 479 := 0;
    variable x_length : integer range 0 to 639 := 0;
  begin
    if (display_en = '1') then
      if (column mod 5 = 0 or row mod 6 = 0) then
        VGA_R <= (others => '1');
        VGA_G <= (others => '0');
        VGA_B <= (others => '0');
      else
        VGA_R <= (others => '0');
        VGA_G <= (others => '0');
        VGA_B <= (others => '1');
      end if;

    else
      VGA_R <= (others => '0');
      VGA_G <= (others => '0');
      VGA_B <= (others => '0');
    end if;
  end process;
  
  vga_adpater_1 : vga_adapter
    port map(
      pixel_clk => clk,
      reset_n => KEY(3),
      h_sync => VGA_HS,
      v_sync => VGA_VS,
      blank_n => VGA_BLANK_N,
      sync_n => VGA_SYNC_N,
      display_en => display_en,
      column => column,
      row => row
    );
END RTL;

